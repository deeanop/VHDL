library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity tb_not_gate is
end tb_not_gate;

architecture test of tb_not_gate is
	signal A, Y : STD_LOGIC;
begin
	uut: entity work.not_gate
		port map (
			A => A,
			Y => Y
		);
	stim_proc: process
	begin
		A <= '0'; wait for 10 ns;
		A <= '1'; wait for 10 ns;
		wait;
	end process;
end test;
	 