library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity not_gate is
	Port (
		A : in STD_LOGIC;
		Y : out STD_LOGIC
	);
end not_gate;

architecture behavior of not_gate is
begin
	Y <= NOT A;
end behavior;
